------------------------------------------------------------------------------------------------------------------------
-- True Dual Port RAM - 32Kb x 1k
------------------------------------------------------------------------------------------------------------------------
--Standard Libraries
library ieee;
use ieee.std_logic_1164.all;
--
Library UNISIM;
use UNISIM.vcomponents.all;

entity true_dualportbe_ram is
    Port (
        --Port A
      rsta_i    : in  std_logic;                        -- 1-bit A port set/reset input
      clka_i    : in  std_logic;                        -- 1-bit A port clock input
      wrena_i   : in  std_logic_vector(3 downto 0);     -- 4-bit A port write enable input
      rdena_i   : in  std_logic;                        -- 1-bit A port enable input
      dataa_i   : in  std_logic_vector(31 downto 0);    -- 32-bit A port data input
      dataa_o   : out std_logic_vector(31 downto 0);    -- 32-bit A port data output
      addra_i   : in  std_logic_vector(9 downto 0);     -- 12-bit A port address input
      --Port B
      rstb_i    : in  std_logic;                        -- 1-bit B port set/reset input
      clkb_i    : in  std_logic;                        -- 1 bit B port clock input
      wrenb_i   : in  std_logic_vector(3 downto 0);     -- 4-bit B port write enable input
      rdenb_i   : in  std_logic;                        -- 1-bit B port enable input
      datab_i   : in  std_logic_vector(31 downto 0);    -- 32-bit B port data input
      datab_o   : out std_logic_vector(31 downto 0);    -- 32-bit B port data output
      addrb_i   : in  std_logic_vector(9 downto 0)      -- 12-bit B port address input
    );

end true_dualportbe_ram;

architecture rtl of true_dualportbe_ram is

  --Optional ports
  --signal CASCADEOUTLATA : std_logic:='0';
  -- 1-bit cascade A latch output
  --signal CASCADEOUTLATB : std_logic:='0';
  -- 1-bit cascade B latch output
  --signal CASCADEOUTREGA : std_logic:='0';
  -- 1-bit cascade A register output
  --signal CASCADEOUTREGB : std_logic:='0';
  -- 1-bit cascade B register output
  signal DOPA           : std_logic_vector(3 downto 0):=(others=>'0');   -- 4-bit A port parity data output
  signal DOPB           : std_logic_vector(3 downto 0):=(others=>'0');   -- 4-bit B port parity data output
  signal CASCADEINLATA  : std_logic:='0';                        -- 1-bit cascade A latch input
  signal CASCADEINLATB  : std_logic:='0';                          -- 1-bit cascade B latch input
  signal CASCADEINREGA  : std_logic:='0';                          -- 1-bit cascade A register input
  signal CASCADEINREGB  : std_logic:='0';                          -- 1-bit cascade B register input
  signal DIPA           : std_logic_vector(3 downto 0):=(others=>'0');            -- 4-bit A port parity data input
  signal DIPB           : std_logic_vector(3 downto 0):=(others=>'0');            -- 4-bit B port parity data input
  signal REGCEA         : std_logic:='0';                          -- 1-bit A port register enable input
  signal REGCEB         : std_logic:='0';                          -- 1-bit B port register enable input
  signal addra_s        : std_logic_vector(15 downto 0);
  signal addrb_s        : std_logic_vector(15 downto 0);
begin


-- ADDR pins must be 16-bits wide. However, valid addresses for non-cascadable block RAM
-- are only found on pin 14 to (15 - address width). The remaining pins, including pin 15, should be tied High.
    addra_s <= '1'&addra_i&"11111";
    addrb_s <= '1'&addrb_i&"11111";

-- RAMB36: 32k+4k Parity Paramatizable True Dual-Port BlockRAM
-- Virtex-5
-- Xilinx HDL Libraries Guide, version 12.4
  RAMB36_inst : RAMB36
  generic map (
    DOA_REG     => 0, -- Optional output register on A port (0 or 1)
    DOB_REG     => 0, -- Optional output register on B port (0 or 1)
    INIT_A      => X"000000000", -- Initial values on A output port
    INIT_B      => X"000000000", -- Initial values on B output port
    RAM_EXTENSION_A  => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
    RAM_EXTENSION_B  => "NONE", -- "UPPER", "LOWER" or "NONE" when cascaded
    READ_WIDTH_A     => 36,
    -- Valid values are 1, 2, 4, 9, 18, or 36
    READ_WIDTH_B     => 36,
    -- Valid values are 1, 2, 4, 9, 18, or 36
    SIM_COLLISION_CHECK   => "ALL", -- Collision check enable "ALL", "WARNING_ONLY",
    -- "GENERATE_X_ONLY" or "NONE"
    SIM_MODE     => "SAFE", -- Simulation: "SAFE" vs "FAST", see "Synthesis and Simulation
    -- Design Guide" for details

    SRVAL_A   => X"000000000",
    -- Set/Reset value for A port output
    SRVAL_B   => X"000000000",
    -- Set/Reset value for B port output
    WRITE_MODE_A   => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    WRITE_MODE_B   => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    WRITE_WIDTH_A  => 36, -- Valid values are 1, 2, 3, 4, 9, 18, 36
    WRITE_WIDTH_B  => 36, -- Valid values are 1, 2, 3, 4, 9, 18, 36
    -- The following INIT_xx declarations specify the initial contents of the RAM
    INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
    -- The next set of INITP_xx are for the parity bits
    INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
  port map (
    --CASCADEOUTLATA   => CASCADEOUTLATA,
    -- 1-bit cascade A latch output
    --CASCADEOUTLATB   => CASCADEOUTLATB,
    -- 1-bit cascade B latch output
    --CASCADEOUTREGA   => CASCADEOUTREGA,
    -- 1-bit cascade A register output
    --CASCADEOUTREGB   => CASCADEOUTREGB,
    -- 1-bit cascade B register output
    DOA     => dataa_o,                 -- 32-bit A port data output
    DOB     => datab_o,                 -- 32-bit B port data output
    DOPA    => DOPA,                    -- 4-bit A port parity data output
    DOPB    => DOPB,                    -- 4-bit B port parity data output
    ADDRA   => addra_s,                 -- 16-bit A port address input
    ADDRB   => addrb_s,                 -- 16-bit B port address input
    CASCADEINLATA   => CASCADEINLATA,   -- 1-bit cascade A latch input
    CASCADEINLATB   => CASCADEINLATB,   -- 1-bit cascade B latch input
    CASCADEINREGA   => CASCADEINREGA,   -- 1-bit cascade A register input
    CASCADEINREGB   => CASCADEINREGB,   -- 1-bit cascade B register input
    CLKA    => clka_i,                  -- 1-bit A port clock input
    CLKB    => clkb_i,                  -- 1 bit B port clock input
    DIA     => dataa_i,                 -- 32-bit A port data input
    DIB     => datab_i,                 -- 32-bit B port data input
    DIPA    => DIPA,                    -- 4-bit A port parity data input
    DIPB    => DIPB,                    -- 4-bit B port parity data input
    ENA     => rdena_i,                 -- 1-bit A port enable input
    ENB     => rdenb_i,                 -- 1-bit B port enable input
    REGCEA  => REGCEA,                  -- 1-bit A port register enable input
    REGCEB  => REGCEB,                  -- 1-bit B port register enable input
    SSRA    => rsta_i,                  -- 1-bit A port set/reset input
    SSRB    => rstb_i,                  -- 1-bit B port set/reset input
    WEA     => wrena_i,                 -- 4-bit A port write enable input
    WEB     => wrenb_i                  -- 4-bit B port write enable input
  );
  -- End of RAMB36_inst instantiation

end rtl;
